package util_pkg;
  
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "timescale.sv"
    `include "config_macro.svh"

endpackage