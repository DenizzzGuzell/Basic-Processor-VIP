package alu_agent_pkg_hdl;

  import util_pkg::*;
  
  `include "timescale.sv"
  `include "alu_macros.svh"

endpackage