package agent_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "./../utils/config_macro.svh"

	`include "./../sequences/sequence_item.svh"
	`include "agent_cfg.svh"
	`include "driver.svh"
	`include "monitor.svh"
	`include "sequencer.svh"
	`include "agent.svh"
	`include "./../sequences/sequence.svh"
endpackage: agent_pkg
