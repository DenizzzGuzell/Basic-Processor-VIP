package alu_agent_pkg;

	import uvm_pkg::*;
	import util_pkg::*;
	`include "uvm_macros.svh"
	`include "config_macro.svh"
	`include "timescale.sv"
	`include "alu_macros.svh"

	`include "alu_sequence_item.svh"
	`include "alu_agent_cfg.svh"
	`include "alu_driver.svh"
	`include "alu_monitor.svh"
	`include "alu_agent.svh"
	`include "./../sequences/alu_base_sequence.svh"
endpackage: alu_agent_pkg
