package alu_test_lib_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"

	import util_pkg::*;
	`include "timescale.sv"

	import alu_env_pkg::*;
	import alu_agent_pkg::*;
	`include "alu_test_base.svh"
	`include "alu_system_test.svh"

endpackage: alu_test_lib_pkg
