`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: YONGATEK
// Engineer:
//
// Create Date: 11/08/2022 11:38:27 AM
// Design Name:
// Module Name: simple_ALU
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module simple_ALU(input i_clk,
				  input i_rst,
				  input logic  [15:0] i_memData,
				  output logic  [15:0]  o_memData,
				  output logic [15:0] o_memAddr,
				  output logic o_memWrEnable);
endmodule
